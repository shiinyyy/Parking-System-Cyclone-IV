module servo (

);
